module Load(in, result);
  input [31:0] in;
  output [31:0] result;
  assign result = in;
endmodule
