`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    07:50:27 11/14/2021 
// Design Name: 
// Module Name:    TopLevelMemoryControl 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module TopLevelMemoryControl(src1,src2,opCode,RW,AddbusDataAcess,
							dataBusIn,dataBusOut,dataOutLDR,PC);
							

endmodule
