module MovReg(in1, result);
  input [31:0] in1;
  output [31:0] result;
  assign result = in1;
endmodule
