module MovN(imvalue, result);
  input [15:0] imvalue;
  output [31:0] result;
  assign result = imvalue;
endmodule
