module 

reg [31:0] machine_code;

// wire ?? ;



initial begin

machineCode = 0;

#5 machineCode = ;
#5 machineCode = ;
#5 machineCode = ;
#5 machineCode = ;
#5 machineCode = ;
#5 machineCode = ;
#5 machineCode = ;
#5 machineCode = ;
#5 machineCode = ;
#5 machineCode = ;
#5 machineCode = ;
#5 machineCode = ;
#5 machineCode = ;
#5 machineCode = ;
#5 machineCode = ;
#5 machineCode = ;
#5 machineCode = ;
#5 machineCode = ;
end
initial begin
    $monitor(,);
end

endmodule
