`timescale 1ns / 1ps
//Condition-OPCode-S-Destination-/Src1/Src2/ShiftROR/3bits/-ShiftRORControl
//4-4-1-4-/4/4/5/3/-3
// 4/4/5/3 Imidiate value 16 bits
module InstructionDecoder();


endmodule
